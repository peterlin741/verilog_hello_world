module hello_world;

  initial begin
    $display("Hello, World!"); // Display the message
    $finish;                  // Terminate the simulation
  end

endmodule